// `timescale 1ns/1ns
package alu_package;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Files
    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "subscriber.sv"
    `include "env.sv"
    `include "test.sv"
endpackage: alu_package